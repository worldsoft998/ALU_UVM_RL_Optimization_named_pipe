package alu_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "alu_seq_item.sv"
  `include "alu_driver.sv"
  `include "alu_monitor.sv"
  `include "alu_sequencer.sv"
  `include "alu_agent.sv"
  `include "alu_scoreboard.sv"
  `include "alu_coverage.sv"
  `include "ai_bridge.sv"
  `include "alu_env.sv"
  `include "alu_base_seq.sv"
  `include "alu_random_seq.sv"
  `include "alu_base_test.sv"
  `include "alu_random_test.sv"
endpackage